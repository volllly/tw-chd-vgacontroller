configuration content_ctrl_cfg of content_ctrl is
  for struc_mem1 
  end for;
end configuration;