configuration content_ctrl_cfg of content_ctrl is
  for rtl_mem2
  end for;
end configuration;