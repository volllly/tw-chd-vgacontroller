configuration vga_controler_top_cfg of vga_controler_top is
  for struc_mem1 
  end for;
end configuration;