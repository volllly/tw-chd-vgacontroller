configuration tb_vga_cfg of tb_vga is
  for sim_mem1 
  end for;
end configuration;